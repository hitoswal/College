---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.LCD_String_DataType.all;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
entity LCD_String is 
Port(	Input : in std_logic_vector(5 downto 0);
		In_Data_N : in std_logic_vector(3 downto 0);
		In_Data_D : in std_logic_vector(3 downto 0);
		In_Data_Q : in std_logic_vector(3 downto 0);
		Output : out character_string);
end LCD_String;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
architecture ckt of LCD_String is
begin
process(Input)
begin
---------------------------------------------------------------------------------
if Input = "000000" then
Output <= (
-- Line 1----MACHINE CLOSED
   X"20",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",
	X"20",X"43",X"4C",X"4F",X"53",X"45",X"44",X"20",
-- Line 2----SWITCH ON SW1
   X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"20",
	X"4F",X"4E",X"20",X"53",X"57",X"31",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "000001" then
Output <= (
-- Line 1----WELCOME!!!
   X"20",X"20",X"20",X"57",X"45",X"4C",X"43",X"4F",
	X"4D",X"45",X"21",X"21",X"21",X"20",X"20",X"20",
-- Line 2----CHIPS:30 COCA:25
   X"43",X"48",X"49",X"50",X"53",X"3A",X"33",X"30",
	X"20",X"43",X"4F",X"43",X"41",X"3A",X"32",X"35");
---------------------------------------------------------------------------------
elsif Input = "000010" then
Output <= (
-- Line 1-----RET N:X D:X Q:X
   X"52",X"45",X"54",X"20",X"4E",X"3A",X"0" & In_Data_N,X"20",X"44",
	X"3A",X"0" & In_Data_D,X"20",X"51",X"3A",X"0" & In_Data_Q,X"20",
-- Line 2----CHIPS:30 COLA:25
   X"43",X"48",X"49",X"50",X"53",X"3A",X"33",X"30",
	X"20",X"43",X"4F",X"43",X"41",X"3A",X"32",X"35");
---------------------------------------------------------------------------------
elsif Input = "000011" then
Output <= (
-- Line 1-----MAX AMOUNT 2.00
   X"4D",X"41",X"58",X"20",X"41",X"4D",X"4F",X"55",
	X"4E",X"54",X"20",X"32",X"2E",X"30",X"30",X"20",
-- Line 2-----SELECT PRODUCT
   X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"50",
	X"52",X"4F",X"44",X"55",X"43",X"54",X"20",X"20");
---------------------------------------------------------------------------------
end if;
end process;
end ckt;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------