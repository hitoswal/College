---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.LCD_String_DataType.all;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
entity LCD_String is 
Port(	Input : in std_logic_vector(3 downto 0);
		In_Data : in std_logic_vector(8 downto 0);
		Output : out character_string);
end LCD_String;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
architecture ckt of LCD_String is
begin
process(Input)
begin
---------------------------------------------------------------------------------
if Input = "0000" then
Output <= (
-- Line 1----SEQ AND INPUT.
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0001" then
Output <= (
-- Line 1----BIT1
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"2D",X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0010" then
Output <= (
-- Line 1-----BIT2
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"2D",X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0011" then
Output <= (
-- Line 1-----BIT3
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"2D",
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0100" then
Output <= (
-- Line 1-----BIT4
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"2D",X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0101" then
Output <= (
-- Line 1-----BIT5
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"2D",X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0110" then
Output <= (
-- Line 1-----BIT6
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"2D",X"0" & "000" & In_Data(2),
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "0111" then
Output <= (
-- Line 1-----BIT7
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"2D",
	X"0" & "000" & In_Data(1),X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "1000" then
Output <= (
-- Line 1-----BIT8
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"49",X"4E",X"3A",X"20",X"0" & "000" & In_Data(8),X"0" & "000" & In_Data(7),X"0" & "000" & In_Data(6),
	X"0" & "000" & In_Data(5),X"0" & "000" & In_Data(4),X"0" & "000" & In_Data(3),X"0" & "000" & In_Data(2),
	X"2D",X"0" & "000" & In_Data(0),X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "1010" then
Output <= (
-- Line 1-----FAIL
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"20",X"20",X"20",X"20", X"20",X"46",X"41",X"49",
	X"4C",X"21",X"21",X"20",X"20",X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "1011" then
Output <= (
-- Line 1-----SUCCESS
   X"53",X"45",X"51",X"3A",X"20",X"31",X"31",X"30",
	X"31",X"31",X"30",X"31",X"30",X"31",X"20",X"20",
-- Line 2
   X"20",X"20",X"20",X"53", X"55",X"43",X"43",X"45",
	X"53",X"53",X"21",X"21",X"21",X"20",X"20",X"20");
---------------------------------------------------------------------------------
end if;
end process;
end ckt;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------