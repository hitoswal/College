---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.LCD_String_DataType.all;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
entity LCD_String is 
Port(	Input : in std_logic_vector(2 downto 0);
		Output : out character_string);
end LCD_String;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------
architecture ckt of LCD_String is
begin
process(Input)
begin
---------------------------------------------------------------------------------
if Input = "000" then
Output <= (
-- Line 1----WELCOME!! PRESS
   X"57",X"45",X"4C",X"43",X"4F",X"4D",X"45",X"21",
	X"21",X"20",X"50",X"52",X"45",X"53",X"53",X"20",
-- Line 2----KEY 3 TO START
   X"4B",X"45",X"59",X"20",X"33",X"20",X"54",X"4F",
	X"20",X"53",X"54",X"41",X"52",X"54",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "001" then
Output <= (
-- Line 1----PRESS KEY 3 TO 
   X"50",X"52",X"45",X"53",X"53",X"20",X"4B",X"45",
	X"59",X"20",X"33",X"20",X"54",X"4F",X"20",X"20",
-- Line 2----STOP
   X"53",X"54",X"4F",X"50",X"20",X"20",X"20",X"20",
	X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "010" then
Output <= (
-- Line 1-----YOU WIN!!
   X"59",X"4F",X"55",X"20",X"57",X"49",X"4E",X"21",
	X"21",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
-- Line 2----
   X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
	X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20");
---------------------------------------------------------------------------------
elsif Input = "011" then
Output <= (
-- Line 1-----YOU LOSE!!
   X"59",X"4F",X"55",X"20",X"4C",X"4F",X"53",X"45",
	X"21",X"21",X"20",X"20",X"20",X"20",X"20",X"20",
-- Line 2-----
   X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
	X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20");
---------------------------------------------------------------------------------
end if;
end process;
end ckt;
---------------------------------------------------------------------------------
---------------------------------------------------------------------------------