/*Name: Hitesh Vijay Oswal and Kausthub Chaudhari*/ 
module FullAdder(
    input A,
    input B,
    input Cin,
    output S
    );

assign S = A ^ B ^ Cin;

endmodule
